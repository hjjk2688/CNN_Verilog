`timescale 1ns / 1ps

// Generated from: train_4.bmp (Scaled by 127)
module image_rom (
    input wire [9:0] addr,
    output reg [7:0] dout
);

    always @(*) begin
        case(addr)
            10'd0: dout = 8'h00;
            10'd1: dout = 8'h00;
            10'd2: dout = 8'h00;
            10'd3: dout = 8'h00;
            10'd4: dout = 8'h00;
            10'd5: dout = 8'h00;
            10'd6: dout = 8'h00;
            10'd7: dout = 8'h00;
            10'd8: dout = 8'h00;
            10'd9: dout = 8'h00;
            10'd10: dout = 8'h00;
            10'd11: dout = 8'h00;
            10'd12: dout = 8'h00;
            10'd13: dout = 8'h00;
            10'd14: dout = 8'h00;
            10'd15: dout = 8'h00;
            10'd16: dout = 8'h00;
            10'd17: dout = 8'h00;
            10'd18: dout = 8'h00;
            10'd19: dout = 8'h00;
            10'd20: dout = 8'h00;
            10'd21: dout = 8'h00;
            10'd22: dout = 8'h00;
            10'd23: dout = 8'h00;
            10'd24: dout = 8'h00;
            10'd25: dout = 8'h00;
            10'd26: dout = 8'h00;
            10'd27: dout = 8'h00;
            10'd28: dout = 8'h00;
            10'd29: dout = 8'h00;
            10'd30: dout = 8'h00;
            10'd31: dout = 8'h00;
            10'd32: dout = 8'h00;
            10'd33: dout = 8'h00;
            10'd34: dout = 8'h00;
            10'd35: dout = 8'h00;
            10'd36: dout = 8'h00;
            10'd37: dout = 8'h00;
            10'd38: dout = 8'h00;
            10'd39: dout = 8'h00;
            10'd40: dout = 8'h00;
            10'd41: dout = 8'h00;
            10'd42: dout = 8'h00;
            10'd43: dout = 8'h00;
            10'd44: dout = 8'h00;
            10'd45: dout = 8'h00;
            10'd46: dout = 8'h00;
            10'd47: dout = 8'h00;
            10'd48: dout = 8'h00;
            10'd49: dout = 8'h00;
            10'd50: dout = 8'h00;
            10'd51: dout = 8'h00;
            10'd52: dout = 8'h00;
            10'd53: dout = 8'h00;
            10'd54: dout = 8'h00;
            10'd55: dout = 8'h00;
            10'd56: dout = 8'h00;
            10'd57: dout = 8'h00;
            10'd58: dout = 8'h00;
            10'd59: dout = 8'h00;
            10'd60: dout = 8'h00;
            10'd61: dout = 8'h00;
            10'd62: dout = 8'h00;
            10'd63: dout = 8'h00;
            10'd64: dout = 8'h00;
            10'd65: dout = 8'h00;
            10'd66: dout = 8'h00;
            10'd67: dout = 8'h00;
            10'd68: dout = 8'h00;
            10'd69: dout = 8'h00;
            10'd70: dout = 8'h00;
            10'd71: dout = 8'h00;
            10'd72: dout = 8'h00;
            10'd73: dout = 8'h00;
            10'd74: dout = 8'h00;
            10'd75: dout = 8'h00;
            10'd76: dout = 8'h00;
            10'd77: dout = 8'h00;
            10'd78: dout = 8'h00;
            10'd79: dout = 8'h00;
            10'd80: dout = 8'h00;
            10'd81: dout = 8'h00;
            10'd82: dout = 8'h00;
            10'd83: dout = 8'h00;
            10'd84: dout = 8'h00;
            10'd85: dout = 8'h00;
            10'd86: dout = 8'h00;
            10'd87: dout = 8'h00;
            10'd88: dout = 8'h00;
            10'd89: dout = 8'h00;
            10'd90: dout = 8'h00;
            10'd91: dout = 8'h00;
            10'd92: dout = 8'h00;
            10'd93: dout = 8'h00;
            10'd94: dout = 8'h00;
            10'd95: dout = 8'h00;
            10'd96: dout = 8'h00;
            10'd97: dout = 8'h00;
            10'd98: dout = 8'h00;
            10'd99: dout = 8'h00;
            10'd100: dout = 8'h00;
            10'd101: dout = 8'h00;
            10'd102: dout = 8'h00;
            10'd103: dout = 8'h00;
            10'd104: dout = 8'h00;
            10'd105: dout = 8'h00;
            10'd106: dout = 8'h00;
            10'd107: dout = 8'h00;
            10'd108: dout = 8'h00;
            10'd109: dout = 8'h00;
            10'd110: dout = 8'h00;
            10'd111: dout = 8'h00;
            10'd112: dout = 8'h00;
            10'd113: dout = 8'h00;
            10'd114: dout = 8'h00;
            10'd115: dout = 8'h00;
            10'd116: dout = 8'h00;
            10'd117: dout = 8'h00;
            10'd118: dout = 8'h00;
            10'd119: dout = 8'h00;
            10'd120: dout = 8'h00;
            10'd121: dout = 8'h00;
            10'd122: dout = 8'h00;
            10'd123: dout = 8'h00;
            10'd124: dout = 8'h00;
            10'd125: dout = 8'h00;
            10'd126: dout = 8'h00;
            10'd127: dout = 8'h00;
            10'd128: dout = 8'h00;
            10'd129: dout = 8'h00;
            10'd130: dout = 8'h00;
            10'd131: dout = 8'h00;
            10'd132: dout = 8'h00;
            10'd133: dout = 8'h00;
            10'd134: dout = 8'h00;
            10'd135: dout = 8'h00;
            10'd136: dout = 8'h00;
            10'd137: dout = 8'h00;
            10'd138: dout = 8'h00;
            10'd139: dout = 8'h00;
            10'd140: dout = 8'h00;
            10'd141: dout = 8'h00;
            10'd142: dout = 8'h00;
            10'd143: dout = 8'h00;
            10'd144: dout = 8'h00;
            10'd145: dout = 8'h00;
            10'd146: dout = 8'h00;
            10'd147: dout = 8'h00;
            10'd148: dout = 8'h00;
            10'd149: dout = 8'h00;
            10'd150: dout = 8'h00;
            10'd151: dout = 8'h00;
            10'd152: dout = 8'h00;
            10'd153: dout = 8'h00;
            10'd154: dout = 8'h00;
            10'd155: dout = 8'h00;
            10'd156: dout = 8'h00;
            10'd157: dout = 8'h00;
            10'd158: dout = 8'h00;
            10'd159: dout = 8'h00;
            10'd160: dout = 8'h00;
            10'd161: dout = 8'h00;
            10'd162: dout = 8'h00;
            10'd163: dout = 8'h00;
            10'd164: dout = 8'h00;
            10'd165: dout = 8'h00;
            10'd166: dout = 8'h00;
            10'd167: dout = 8'h00;
            10'd168: dout = 8'h00;
            10'd169: dout = 8'h00;
            10'd170: dout = 8'h00;
            10'd171: dout = 8'h00;
            10'd172: dout = 8'h00;
            10'd173: dout = 8'h00;
            10'd174: dout = 8'h00;
            10'd175: dout = 8'h00;
            10'd176: dout = 8'h00;
            10'd177: dout = 8'h00;
            10'd178: dout = 8'h00;
            10'd179: dout = 8'h00;
            10'd180: dout = 8'h00;
            10'd181: dout = 8'h00;
            10'd182: dout = 8'h00;
            10'd183: dout = 8'h00;
            10'd184: dout = 8'h00;
            10'd185: dout = 8'h00;
            10'd186: dout = 8'h00;
            10'd187: dout = 8'h00;
            10'd188: dout = 8'h00;
            10'd189: dout = 8'h00;
            10'd190: dout = 8'h00;
            10'd191: dout = 8'h00;
            10'd192: dout = 8'h00;
            10'd193: dout = 8'h00;
            10'd194: dout = 8'h00;
            10'd195: dout = 8'h00;
            10'd196: dout = 8'h00;
            10'd197: dout = 8'h00;
            10'd198: dout = 8'h00;
            10'd199: dout = 8'h00;
            10'd200: dout = 8'h00;
            10'd201: dout = 8'h00;
            10'd202: dout = 8'h00;
            10'd203: dout = 8'h00;
            10'd204: dout = 8'h00;
            10'd205: dout = 8'h00;
            10'd206: dout = 8'h00;
            10'd207: dout = 8'h00;
            10'd208: dout = 8'h1b;
            10'd209: dout = 8'h4a;
            10'd210: dout = 8'h69;
            10'd211: dout = 8'h7e;
            10'd212: dout = 8'h7e;
            10'd213: dout = 8'h38;
            10'd214: dout = 8'h2b;
            10'd215: dout = 8'h4a;
            10'd216: dout = 8'h1b;
            10'd217: dout = 8'h00;
            10'd218: dout = 8'h00;
            10'd219: dout = 8'h00;
            10'd220: dout = 8'h00;
            10'd221: dout = 8'h00;
            10'd222: dout = 8'h00;
            10'd223: dout = 8'h00;
            10'd224: dout = 8'h00;
            10'd225: dout = 8'h00;
            10'd226: dout = 8'h00;
            10'd227: dout = 8'h00;
            10'd228: dout = 8'h00;
            10'd229: dout = 8'h00;
            10'd230: dout = 8'h00;
            10'd231: dout = 8'h00;
            10'd232: dout = 8'h00;
            10'd233: dout = 8'h00;
            10'd234: dout = 8'h00;
            10'd235: dout = 8'h2b;
            10'd236: dout = 8'h74;
            10'd237: dout = 8'h7e;
            10'd238: dout = 8'h7e;
            10'd239: dout = 8'h5e;
            10'd240: dout = 8'h69;
            10'd241: dout = 8'h7e;
            10'd242: dout = 8'h7e;
            10'd243: dout = 8'h7e;
            10'd244: dout = 8'h54;
            10'd245: dout = 8'h00;
            10'd246: dout = 8'h00;
            10'd247: dout = 8'h00;
            10'd248: dout = 8'h00;
            10'd249: dout = 8'h00;
            10'd250: dout = 8'h00;
            10'd251: dout = 8'h00;
            10'd252: dout = 8'h00;
            10'd253: dout = 8'h00;
            10'd254: dout = 8'h00;
            10'd255: dout = 8'h00;
            10'd256: dout = 8'h00;
            10'd257: dout = 8'h00;
            10'd258: dout = 8'h00;
            10'd259: dout = 8'h00;
            10'd260: dout = 8'h00;
            10'd261: dout = 8'h02;
            10'd262: dout = 8'h1c;
            10'd263: dout = 8'h79;
            10'd264: dout = 8'h7e;
            10'd265: dout = 8'h5f;
            10'd266: dout = 8'h20;
            10'd267: dout = 8'h02;
            10'd268: dout = 8'h06;
            10'd269: dout = 8'h5b;
            10'd270: dout = 8'h7e;
            10'd271: dout = 8'h7e;
            10'd272: dout = 8'h3a;
            10'd273: dout = 8'h00;
            10'd274: dout = 8'h00;
            10'd275: dout = 8'h00;
            10'd276: dout = 8'h00;
            10'd277: dout = 8'h00;
            10'd278: dout = 8'h00;
            10'd279: dout = 8'h00;
            10'd280: dout = 8'h00;
            10'd281: dout = 8'h00;
            10'd282: dout = 8'h00;
            10'd283: dout = 8'h00;
            10'd284: dout = 8'h00;
            10'd285: dout = 8'h00;
            10'd286: dout = 8'h00;
            10'd287: dout = 8'h00;
            10'd288: dout = 8'h00;
            10'd289: dout = 8'h30;
            10'd290: dout = 8'h7e;
            10'd291: dout = 8'h7e;
            10'd292: dout = 8'h5b;
            10'd293: dout = 8'h07;
            10'd294: dout = 8'h00;
            10'd295: dout = 8'h00;
            10'd296: dout = 8'h2e;
            10'd297: dout = 8'h7e;
            10'd298: dout = 8'h7e;
            10'd299: dout = 8'h70;
            10'd300: dout = 8'h0a;
            10'd301: dout = 8'h00;
            10'd302: dout = 8'h00;
            10'd303: dout = 8'h00;
            10'd304: dout = 8'h00;
            10'd305: dout = 8'h00;
            10'd306: dout = 8'h00;
            10'd307: dout = 8'h00;
            10'd308: dout = 8'h00;
            10'd309: dout = 8'h00;
            10'd310: dout = 8'h00;
            10'd311: dout = 8'h00;
            10'd312: dout = 8'h00;
            10'd313: dout = 8'h00;
            10'd314: dout = 8'h00;
            10'd315: dout = 8'h00;
            10'd316: dout = 8'h42;
            10'd317: dout = 8'h7e;
            10'd318: dout = 8'h7e;
            10'd319: dout = 8'h49;
            10'd320: dout = 8'h07;
            10'd321: dout = 8'h00;
            10'd322: dout = 8'h00;
            10'd323: dout = 8'h00;
            10'd324: dout = 8'h6b;
            10'd325: dout = 8'h7e;
            10'd326: dout = 8'h7e;
            10'd327: dout = 8'h27;
            10'd328: dout = 8'h00;
            10'd329: dout = 8'h00;
            10'd330: dout = 8'h00;
            10'd331: dout = 8'h00;
            10'd332: dout = 8'h00;
            10'd333: dout = 8'h00;
            10'd334: dout = 8'h00;
            10'd335: dout = 8'h00;
            10'd336: dout = 8'h00;
            10'd337: dout = 8'h00;
            10'd338: dout = 8'h00;
            10'd339: dout = 8'h00;
            10'd340: dout = 8'h00;
            10'd341: dout = 8'h00;
            10'd342: dout = 8'h00;
            10'd343: dout = 8'h3f;
            10'd344: dout = 8'h7e;
            10'd345: dout = 8'h7b;
            10'd346: dout = 8'h58;
            10'd347: dout = 8'h04;
            10'd348: dout = 8'h00;
            10'd349: dout = 8'h00;
            10'd350: dout = 8'h04;
            10'd351: dout = 8'h27;
            10'd352: dout = 8'h7a;
            10'd353: dout = 8'h7e;
            10'd354: dout = 8'h40;
            10'd355: dout = 8'h00;
            10'd356: dout = 8'h00;
            10'd357: dout = 8'h00;
            10'd358: dout = 8'h00;
            10'd359: dout = 8'h00;
            10'd360: dout = 8'h00;
            10'd361: dout = 8'h00;
            10'd362: dout = 8'h00;
            10'd363: dout = 8'h00;
            10'd364: dout = 8'h00;
            10'd365: dout = 8'h00;
            10'd366: dout = 8'h00;
            10'd367: dout = 8'h00;
            10'd368: dout = 8'h00;
            10'd369: dout = 8'h00;
            10'd370: dout = 8'h08;
            10'd371: dout = 8'h74;
            10'd372: dout = 8'h7e;
            10'd373: dout = 8'h58;
            10'd374: dout = 8'h00;
            10'd375: dout = 8'h00;
            10'd376: dout = 8'h00;
            10'd377: dout = 8'h12;
            10'd378: dout = 8'h64;
            10'd379: dout = 8'h7e;
            10'd380: dout = 8'h7e;
            10'd381: dout = 8'h54;
            10'd382: dout = 8'h05;
            10'd383: dout = 8'h00;
            10'd384: dout = 8'h00;
            10'd385: dout = 8'h00;
            10'd386: dout = 8'h00;
            10'd387: dout = 8'h00;
            10'd388: dout = 8'h00;
            10'd389: dout = 8'h00;
            10'd390: dout = 8'h00;
            10'd391: dout = 8'h00;
            10'd392: dout = 8'h00;
            10'd393: dout = 8'h00;
            10'd394: dout = 8'h00;
            10'd395: dout = 8'h00;
            10'd396: dout = 8'h00;
            10'd397: dout = 8'h00;
            10'd398: dout = 8'h0b;
            10'd399: dout = 8'h7e;
            10'd400: dout = 8'h7e;
            10'd401: dout = 8'h0f;
            10'd402: dout = 8'h0b;
            10'd403: dout = 8'h3b;
            10'd404: dout = 8'h62;
            10'd405: dout = 8'h78;
            10'd406: dout = 8'h7e;
            10'd407: dout = 8'h7e;
            10'd408: dout = 8'h7d;
            10'd409: dout = 8'h26;
            10'd410: dout = 8'h00;
            10'd411: dout = 8'h00;
            10'd412: dout = 8'h00;
            10'd413: dout = 8'h00;
            10'd414: dout = 8'h00;
            10'd415: dout = 8'h00;
            10'd416: dout = 8'h00;
            10'd417: dout = 8'h00;
            10'd418: dout = 8'h00;
            10'd419: dout = 8'h00;
            10'd420: dout = 8'h00;
            10'd421: dout = 8'h00;
            10'd422: dout = 8'h00;
            10'd423: dout = 8'h00;
            10'd424: dout = 8'h00;
            10'd425: dout = 8'h00;
            10'd426: dout = 8'h08;
            10'd427: dout = 8'h73;
            10'd428: dout = 8'h7e;
            10'd429: dout = 8'h7e;
            10'd430: dout = 8'h7e;
            10'd431: dout = 8'h7e;
            10'd432: dout = 8'h7e;
            10'd433: dout = 8'h71;
            10'd434: dout = 8'h71;
            10'd435: dout = 8'h7e;
            10'd436: dout = 8'h73;
            10'd437: dout = 8'h00;
            10'd438: dout = 8'h00;
            10'd439: dout = 8'h00;
            10'd440: dout = 8'h00;
            10'd441: dout = 8'h00;
            10'd442: dout = 8'h00;
            10'd443: dout = 8'h00;
            10'd444: dout = 8'h00;
            10'd445: dout = 8'h00;
            10'd446: dout = 8'h00;
            10'd447: dout = 8'h00;
            10'd448: dout = 8'h00;
            10'd449: dout = 8'h00;
            10'd450: dout = 8'h00;
            10'd451: dout = 8'h00;
            10'd452: dout = 8'h00;
            10'd453: dout = 8'h00;
            10'd454: dout = 8'h00;
            10'd455: dout = 8'h1b;
            10'd456: dout = 8'h75;
            10'd457: dout = 8'h7e;
            10'd458: dout = 8'h6c;
            10'd459: dout = 8'h45;
            10'd460: dout = 8'h15;
            10'd461: dout = 8'h0c;
            10'd462: dout = 8'h60;
            10'd463: dout = 8'h7e;
            10'd464: dout = 8'h47;
            10'd465: dout = 8'h00;
            10'd466: dout = 8'h00;
            10'd467: dout = 8'h00;
            10'd468: dout = 8'h00;
            10'd469: dout = 8'h00;
            10'd470: dout = 8'h00;
            10'd471: dout = 8'h00;
            10'd472: dout = 8'h00;
            10'd473: dout = 8'h00;
            10'd474: dout = 8'h00;
            10'd475: dout = 8'h00;
            10'd476: dout = 8'h00;
            10'd477: dout = 8'h00;
            10'd478: dout = 8'h00;
            10'd479: dout = 8'h00;
            10'd480: dout = 8'h00;
            10'd481: dout = 8'h00;
            10'd482: dout = 8'h00;
            10'd483: dout = 8'h00;
            10'd484: dout = 8'h00;
            10'd485: dout = 8'h00;
            10'd486: dout = 8'h00;
            10'd487: dout = 8'h00;
            10'd488: dout = 8'h00;
            10'd489: dout = 8'h1f;
            10'd490: dout = 8'h7f;
            10'd491: dout = 8'h7e;
            10'd492: dout = 8'h36;
            10'd493: dout = 8'h00;
            10'd494: dout = 8'h00;
            10'd495: dout = 8'h00;
            10'd496: dout = 8'h00;
            10'd497: dout = 8'h00;
            10'd498: dout = 8'h00;
            10'd499: dout = 8'h00;
            10'd500: dout = 8'h00;
            10'd501: dout = 8'h00;
            10'd502: dout = 8'h00;
            10'd503: dout = 8'h00;
            10'd504: dout = 8'h00;
            10'd505: dout = 8'h00;
            10'd506: dout = 8'h00;
            10'd507: dout = 8'h00;
            10'd508: dout = 8'h00;
            10'd509: dout = 8'h00;
            10'd510: dout = 8'h00;
            10'd511: dout = 8'h00;
            10'd512: dout = 8'h00;
            10'd513: dout = 8'h00;
            10'd514: dout = 8'h00;
            10'd515: dout = 8'h00;
            10'd516: dout = 8'h00;
            10'd517: dout = 8'h23;
            10'd518: dout = 8'h7e;
            10'd519: dout = 8'h7e;
            10'd520: dout = 8'h0a;
            10'd521: dout = 8'h00;
            10'd522: dout = 8'h00;
            10'd523: dout = 8'h00;
            10'd524: dout = 8'h00;
            10'd525: dout = 8'h00;
            10'd526: dout = 8'h00;
            10'd527: dout = 8'h00;
            10'd528: dout = 8'h00;
            10'd529: dout = 8'h00;
            10'd530: dout = 8'h00;
            10'd531: dout = 8'h00;
            10'd532: dout = 8'h00;
            10'd533: dout = 8'h00;
            10'd534: dout = 8'h00;
            10'd535: dout = 8'h00;
            10'd536: dout = 8'h00;
            10'd537: dout = 8'h00;
            10'd538: dout = 8'h00;
            10'd539: dout = 8'h00;
            10'd540: dout = 8'h00;
            10'd541: dout = 8'h00;
            10'd542: dout = 8'h00;
            10'd543: dout = 8'h00;
            10'd544: dout = 8'h00;
            10'd545: dout = 8'h00;
            10'd546: dout = 8'h7e;
            10'd547: dout = 8'h7e;
            10'd548: dout = 8'h0a;
            10'd549: dout = 8'h00;
            10'd550: dout = 8'h00;
            10'd551: dout = 8'h00;
            10'd552: dout = 8'h00;
            10'd553: dout = 8'h00;
            10'd554: dout = 8'h00;
            10'd555: dout = 8'h00;
            10'd556: dout = 8'h00;
            10'd557: dout = 8'h00;
            10'd558: dout = 8'h00;
            10'd559: dout = 8'h00;
            10'd560: dout = 8'h00;
            10'd561: dout = 8'h00;
            10'd562: dout = 8'h00;
            10'd563: dout = 8'h00;
            10'd564: dout = 8'h00;
            10'd565: dout = 8'h00;
            10'd566: dout = 8'h00;
            10'd567: dout = 8'h00;
            10'd568: dout = 8'h00;
            10'd569: dout = 8'h00;
            10'd570: dout = 8'h00;
            10'd571: dout = 8'h00;
            10'd572: dout = 8'h00;
            10'd573: dout = 8'h23;
            10'd574: dout = 8'h7e;
            10'd575: dout = 8'h7e;
            10'd576: dout = 8'h0a;
            10'd577: dout = 8'h00;
            10'd578: dout = 8'h00;
            10'd579: dout = 8'h00;
            10'd580: dout = 8'h00;
            10'd581: dout = 8'h00;
            10'd582: dout = 8'h00;
            10'd583: dout = 8'h00;
            10'd584: dout = 8'h00;
            10'd585: dout = 8'h00;
            10'd586: dout = 8'h00;
            10'd587: dout = 8'h00;
            10'd588: dout = 8'h00;
            10'd589: dout = 8'h00;
            10'd590: dout = 8'h00;
            10'd591: dout = 8'h00;
            10'd592: dout = 8'h00;
            10'd593: dout = 8'h00;
            10'd594: dout = 8'h00;
            10'd595: dout = 8'h00;
            10'd596: dout = 8'h00;
            10'd597: dout = 8'h00;
            10'd598: dout = 8'h00;
            10'd599: dout = 8'h00;
            10'd600: dout = 8'h00;
            10'd601: dout = 8'h35;
            10'd602: dout = 8'h7e;
            10'd603: dout = 8'h7e;
            10'd604: dout = 8'h0a;
            10'd605: dout = 8'h00;
            10'd606: dout = 8'h00;
            10'd607: dout = 8'h00;
            10'd608: dout = 8'h00;
            10'd609: dout = 8'h00;
            10'd610: dout = 8'h00;
            10'd611: dout = 8'h00;
            10'd612: dout = 8'h00;
            10'd613: dout = 8'h00;
            10'd614: dout = 8'h00;
            10'd615: dout = 8'h00;
            10'd616: dout = 8'h00;
            10'd617: dout = 8'h00;
            10'd618: dout = 8'h00;
            10'd619: dout = 8'h00;
            10'd620: dout = 8'h00;
            10'd621: dout = 8'h00;
            10'd622: dout = 8'h00;
            10'd623: dout = 8'h00;
            10'd624: dout = 8'h00;
            10'd625: dout = 8'h00;
            10'd626: dout = 8'h00;
            10'd627: dout = 8'h00;
            10'd628: dout = 8'h00;
            10'd629: dout = 8'h16;
            10'd630: dout = 8'h7f;
            10'd631: dout = 8'h7e;
            10'd632: dout = 8'h0a;
            10'd633: dout = 8'h00;
            10'd634: dout = 8'h00;
            10'd635: dout = 8'h00;
            10'd636: dout = 8'h00;
            10'd637: dout = 8'h00;
            10'd638: dout = 8'h00;
            10'd639: dout = 8'h00;
            10'd640: dout = 8'h00;
            10'd641: dout = 8'h00;
            10'd642: dout = 8'h00;
            10'd643: dout = 8'h00;
            10'd644: dout = 8'h00;
            10'd645: dout = 8'h00;
            10'd646: dout = 8'h00;
            10'd647: dout = 8'h00;
            10'd648: dout = 8'h00;
            10'd649: dout = 8'h00;
            10'd650: dout = 8'h00;
            10'd651: dout = 8'h00;
            10'd652: dout = 8'h00;
            10'd653: dout = 8'h00;
            10'd654: dout = 8'h00;
            10'd655: dout = 8'h00;
            10'd656: dout = 8'h00;
            10'd657: dout = 8'h00;
            10'd658: dout = 8'h6d;
            10'd659: dout = 8'h7e;
            10'd660: dout = 8'h1c;
            10'd661: dout = 8'h00;
            10'd662: dout = 8'h00;
            10'd663: dout = 8'h00;
            10'd664: dout = 8'h00;
            10'd665: dout = 8'h00;
            10'd666: dout = 8'h00;
            10'd667: dout = 8'h00;
            10'd668: dout = 8'h00;
            10'd669: dout = 8'h00;
            10'd670: dout = 8'h00;
            10'd671: dout = 8'h00;
            10'd672: dout = 8'h00;
            10'd673: dout = 8'h00;
            10'd674: dout = 8'h00;
            10'd675: dout = 8'h00;
            10'd676: dout = 8'h00;
            10'd677: dout = 8'h00;
            10'd678: dout = 8'h00;
            10'd679: dout = 8'h00;
            10'd680: dout = 8'h00;
            10'd681: dout = 8'h00;
            10'd682: dout = 8'h00;
            10'd683: dout = 8'h00;
            10'd684: dout = 8'h00;
            10'd685: dout = 8'h00;
            10'd686: dout = 8'h30;
            10'd687: dout = 8'h7e;
            10'd688: dout = 8'h5e;
            10'd689: dout = 8'h15;
            10'd690: dout = 8'h00;
            10'd691: dout = 8'h00;
            10'd692: dout = 8'h00;
            10'd693: dout = 8'h00;
            10'd694: dout = 8'h00;
            10'd695: dout = 8'h00;
            10'd696: dout = 8'h00;
            10'd697: dout = 8'h00;
            10'd698: dout = 8'h00;
            10'd699: dout = 8'h00;
            10'd700: dout = 8'h00;
            10'd701: dout = 8'h00;
            10'd702: dout = 8'h00;
            10'd703: dout = 8'h00;
            10'd704: dout = 8'h00;
            10'd705: dout = 8'h00;
            10'd706: dout = 8'h00;
            10'd707: dout = 8'h00;
            10'd708: dout = 8'h00;
            10'd709: dout = 8'h00;
            10'd710: dout = 8'h00;
            10'd711: dout = 8'h00;
            10'd712: dout = 8'h00;
            10'd713: dout = 8'h00;
            10'd714: dout = 8'h07;
            10'd715: dout = 8'h5c;
            10'd716: dout = 8'h7e;
            10'd717: dout = 8'h55;
            10'd718: dout = 8'h05;
            10'd719: dout = 8'h00;
            10'd720: dout = 8'h00;
            10'd721: dout = 8'h00;
            10'd722: dout = 8'h00;
            10'd723: dout = 8'h00;
            10'd724: dout = 8'h00;
            10'd725: dout = 8'h00;
            10'd726: dout = 8'h00;
            10'd727: dout = 8'h00;
            10'd728: dout = 8'h00;
            10'd729: dout = 8'h00;
            10'd730: dout = 8'h00;
            10'd731: dout = 8'h00;
            10'd732: dout = 8'h00;
            10'd733: dout = 8'h00;
            10'd734: dout = 8'h00;
            10'd735: dout = 8'h00;
            10'd736: dout = 8'h00;
            10'd737: dout = 8'h00;
            10'd738: dout = 8'h00;
            10'd739: dout = 8'h00;
            10'd740: dout = 8'h00;
            10'd741: dout = 8'h00;
            10'd742: dout = 8'h00;
            10'd743: dout = 8'h07;
            10'd744: dout = 8'h49;
            10'd745: dout = 8'h7e;
            10'd746: dout = 8'h15;
            10'd747: dout = 8'h00;
            10'd748: dout = 8'h00;
            10'd749: dout = 8'h00;
            10'd750: dout = 8'h00;
            10'd751: dout = 8'h00;
            10'd752: dout = 8'h00;
            10'd753: dout = 8'h00;
            10'd754: dout = 8'h00;
            10'd755: dout = 8'h00;
            10'd756: dout = 8'h00;
            10'd757: dout = 8'h00;
            10'd758: dout = 8'h00;
            10'd759: dout = 8'h00;
            10'd760: dout = 8'h00;
            10'd761: dout = 8'h00;
            10'd762: dout = 8'h00;
            10'd763: dout = 8'h00;
            10'd764: dout = 8'h00;
            10'd765: dout = 8'h00;
            10'd766: dout = 8'h00;
            10'd767: dout = 8'h00;
            10'd768: dout = 8'h00;
            10'd769: dout = 8'h00;
            10'd770: dout = 8'h00;
            10'd771: dout = 8'h00;
            10'd772: dout = 8'h00;
            10'd773: dout = 8'h00;
            10'd774: dout = 8'h00;
            10'd775: dout = 8'h00;
            10'd776: dout = 8'h00;
            10'd777: dout = 8'h00;
            10'd778: dout = 8'h00;
            10'd779: dout = 8'h00;
            10'd780: dout = 8'h00;
            10'd781: dout = 8'h00;
            10'd782: dout = 8'h00;
            10'd783: dout = 8'h00;
            default: dout = 8'h00;
        endcase
    end

endmodule